module sirv_gnrl_buffs (
    
);

endmodule //sirv_gnrl_buffs